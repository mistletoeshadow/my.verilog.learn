`timescale 1ns/1ps

module dds_wave (
    input []
);

endmodule //dds_wave