`timescale 1ns/1ps

module dds_wave (
    input f_clk,
    input rst_n,
    input reg [31:0] f_word,
    input reg [10:0] p_word
    
);



endmodule //dds_wave