library verilog;
use verilog.vl_types.all;
entity dds_tb is
end dds_tb;
