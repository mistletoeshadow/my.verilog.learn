`timescale 1ns/1ps

module dds_wave (
    input [31:0] K,
    input clk,
    input rst_n
);

endmodule //dds_wave