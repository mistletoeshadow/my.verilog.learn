`timescale 1ns/1ps

module dds_wave (
    input [31:0] K,
    input []
);

endmodule //dds_wave