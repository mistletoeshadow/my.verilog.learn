`timescale 1ns/1ps

module dds_wave (
    
);

endmodule //dds_wave