`timescale 1ns/1ps

module dds_wave (
    input [31:0] K,
    input clk
);

endmodule //dds_wave